library verilog;
use verilog.vl_types.all;
entity Divider_vlg_check_tst is
    port(
        overflow        : in     vl_logic;
        Q0              : in     vl_logic;
        Q1              : in     vl_logic;
        Q2              : in     vl_logic;
        Q3              : in     vl_logic;
        Q4              : in     vl_logic;
        Q5              : in     vl_logic;
        Q6              : in     vl_logic;
        Q7              : in     vl_logic;
        Q8              : in     vl_logic;
        Q9              : in     vl_logic;
        Q10             : in     vl_logic;
        Q11             : in     vl_logic;
        Q12             : in     vl_logic;
        Q13             : in     vl_logic;
        Q14             : in     vl_logic;
        Q15             : in     vl_logic;
        Q16             : in     vl_logic;
        Q17             : in     vl_logic;
        Q18             : in     vl_logic;
        Q19             : in     vl_logic;
        Q20             : in     vl_logic;
        Q21             : in     vl_logic;
        Q22             : in     vl_logic;
        Q23             : in     vl_logic;
        S47             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Divider_vlg_check_tst;
