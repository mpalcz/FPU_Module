library verilog;
use verilog.vl_types.all;
entity Divider_vlg_vec_tst is
end Divider_vlg_vec_tst;
