library verilog;
use verilog.vl_types.all;
entity Normalizer_vlg_vec_tst is
end Normalizer_vlg_vec_tst;
