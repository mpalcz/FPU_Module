library verilog;
use verilog.vl_types.all;
entity Divider_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        D4              : in     vl_logic;
        D5              : in     vl_logic;
        D6              : in     vl_logic;
        D7              : in     vl_logic;
        D8              : in     vl_logic;
        D9              : in     vl_logic;
        D10             : in     vl_logic;
        D11             : in     vl_logic;
        D12             : in     vl_logic;
        D13             : in     vl_logic;
        D14             : in     vl_logic;
        D15             : in     vl_logic;
        D16             : in     vl_logic;
        D17             : in     vl_logic;
        D18             : in     vl_logic;
        D19             : in     vl_logic;
        D20             : in     vl_logic;
        D21             : in     vl_logic;
        D22             : in     vl_logic;
        D23             : in     vl_logic;
        R0              : in     vl_logic;
        R1              : in     vl_logic;
        R2              : in     vl_logic;
        R3              : in     vl_logic;
        R4              : in     vl_logic;
        R5              : in     vl_logic;
        R6              : in     vl_logic;
        R7              : in     vl_logic;
        R8              : in     vl_logic;
        R9              : in     vl_logic;
        R10             : in     vl_logic;
        R11             : in     vl_logic;
        R12             : in     vl_logic;
        R13             : in     vl_logic;
        R14             : in     vl_logic;
        R15             : in     vl_logic;
        R16             : in     vl_logic;
        R17             : in     vl_logic;
        R18             : in     vl_logic;
        R19             : in     vl_logic;
        R20             : in     vl_logic;
        R21             : in     vl_logic;
        R22             : in     vl_logic;
        R23             : in     vl_logic;
        Sel             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Divider_vlg_sample_tst;
