library verilog;
use verilog.vl_types.all;
entity Normalizer_vlg_check_tst is
    port(
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        B3              : in     vl_logic;
        B4              : in     vl_logic;
        B5              : in     vl_logic;
        B6              : in     vl_logic;
        B7              : in     vl_logic;
        B8              : in     vl_logic;
        B9              : in     vl_logic;
        B10             : in     vl_logic;
        B11             : in     vl_logic;
        B12             : in     vl_logic;
        B13             : in     vl_logic;
        B14             : in     vl_logic;
        B15             : in     vl_logic;
        B16             : in     vl_logic;
        B17             : in     vl_logic;
        B18             : in     vl_logic;
        B19             : in     vl_logic;
        B20             : in     vl_logic;
        B21             : in     vl_logic;
        B22             : in     vl_logic;
        E0              : in     vl_logic;
        E1              : in     vl_logic;
        E2              : in     vl_logic;
        E3              : in     vl_logic;
        E4              : in     vl_logic;
        E5              : in     vl_logic;
        E6              : in     vl_logic;
        E7              : in     vl_logic;
        Overflow        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Normalizer_vlg_check_tst;
