library verilog;
use verilog.vl_types.all;
entity Multiplier_vlg_sample_tst is
    port(
        Clk             : in     vl_logic;
        En              : in     vl_logic;
        L0              : in     vl_logic;
        L1              : in     vl_logic;
        L2              : in     vl_logic;
        L3              : in     vl_logic;
        L4              : in     vl_logic;
        L5              : in     vl_logic;
        L6              : in     vl_logic;
        L7              : in     vl_logic;
        L8              : in     vl_logic;
        L9              : in     vl_logic;
        L10             : in     vl_logic;
        L11             : in     vl_logic;
        L12             : in     vl_logic;
        L13             : in     vl_logic;
        L14             : in     vl_logic;
        L15             : in     vl_logic;
        L16             : in     vl_logic;
        L17             : in     vl_logic;
        L18             : in     vl_logic;
        L19             : in     vl_logic;
        L20             : in     vl_logic;
        L21             : in     vl_logic;
        L22             : in     vl_logic;
        L23             : in     vl_logic;
        Multiplicand0   : in     vl_logic;
        Multiplicand1   : in     vl_logic;
        Multiplicand2   : in     vl_logic;
        Multiplicand3   : in     vl_logic;
        Multiplicand4   : in     vl_logic;
        Multiplicand5   : in     vl_logic;
        Multiplicand6   : in     vl_logic;
        Multiplicand7   : in     vl_logic;
        Multiplicand8   : in     vl_logic;
        Multiplicand9   : in     vl_logic;
        Multiplicand10  : in     vl_logic;
        Multiplicand11  : in     vl_logic;
        Multiplicand12  : in     vl_logic;
        Multiplicand13  : in     vl_logic;
        Multiplicand14  : in     vl_logic;
        Multiplicand15  : in     vl_logic;
        Multiplicand16  : in     vl_logic;
        Multiplicand17  : in     vl_logic;
        Multiplicand18  : in     vl_logic;
        Multiplicand19  : in     vl_logic;
        Multiplicand20  : in     vl_logic;
        Multiplicand21  : in     vl_logic;
        Multiplicand22  : in     vl_logic;
        Multiplicand23  : in     vl_logic;
        Sel             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Multiplier_vlg_sample_tst;
