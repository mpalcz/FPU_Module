library verilog;
use verilog.vl_types.all;
entity Divider is
    port(
        Q22             : out    vl_logic;
        Q0              : out    vl_logic;
        clk             : in     vl_logic;
        S47             : out    vl_logic;
        R0              : in     vl_logic;
        Sel             : in     vl_logic;
        R1              : in     vl_logic;
        R2              : in     vl_logic;
        R3              : in     vl_logic;
        R4              : in     vl_logic;
        R5              : in     vl_logic;
        R6              : in     vl_logic;
        R7              : in     vl_logic;
        R8              : in     vl_logic;
        R9              : in     vl_logic;
        R10             : in     vl_logic;
        R11             : in     vl_logic;
        R12             : in     vl_logic;
        R13             : in     vl_logic;
        R14             : in     vl_logic;
        R15             : in     vl_logic;
        R16             : in     vl_logic;
        R17             : in     vl_logic;
        R18             : in     vl_logic;
        R19             : in     vl_logic;
        R20             : in     vl_logic;
        R21             : in     vl_logic;
        R22             : in     vl_logic;
        R23             : in     vl_logic;
        D23             : in     vl_logic;
        D22             : in     vl_logic;
        D21             : in     vl_logic;
        D20             : in     vl_logic;
        D19             : in     vl_logic;
        D18             : in     vl_logic;
        D17             : in     vl_logic;
        D16             : in     vl_logic;
        D15             : in     vl_logic;
        D14             : in     vl_logic;
        D13             : in     vl_logic;
        D12             : in     vl_logic;
        D11             : in     vl_logic;
        D10             : in     vl_logic;
        D9              : in     vl_logic;
        D8              : in     vl_logic;
        D7              : in     vl_logic;
        D6              : in     vl_logic;
        D5              : in     vl_logic;
        D4              : in     vl_logic;
        D3              : in     vl_logic;
        D2              : in     vl_logic;
        D1              : in     vl_logic;
        D0              : in     vl_logic;
        Q21             : out    vl_logic;
        Q20             : out    vl_logic;
        Q19             : out    vl_logic;
        Q18             : out    vl_logic;
        Q17             : out    vl_logic;
        Q16             : out    vl_logic;
        Q15             : out    vl_logic;
        Q14             : out    vl_logic;
        Q13             : out    vl_logic;
        Q12             : out    vl_logic;
        Q11             : out    vl_logic;
        Q10             : out    vl_logic;
        Q9              : out    vl_logic;
        Q8              : out    vl_logic;
        Q7              : out    vl_logic;
        Q6              : out    vl_logic;
        Q5              : out    vl_logic;
        Q4              : out    vl_logic;
        Q3              : out    vl_logic;
        Q2              : out    vl_logic;
        Q1              : out    vl_logic;
        Q23             : out    vl_logic;
        overflow        : out    vl_logic
    );
end Divider;
