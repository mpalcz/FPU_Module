library verilog;
use verilog.vl_types.all;
entity Multiplier_vlg_check_tst is
    port(
        bit_out         : in     vl_logic;
        mux0            : in     vl_logic;
        mux1            : in     vl_logic;
        mux2            : in     vl_logic;
        mux3            : in     vl_logic;
        mux4            : in     vl_logic;
        mux5            : in     vl_logic;
        mux6            : in     vl_logic;
        mux7            : in     vl_logic;
        Overflow        : in     vl_logic;
        prod0           : in     vl_logic;
        prod1           : in     vl_logic;
        prod2           : in     vl_logic;
        prod3           : in     vl_logic;
        prod4           : in     vl_logic;
        prod5           : in     vl_logic;
        prod6           : in     vl_logic;
        prod7           : in     vl_logic;
        prod8           : in     vl_logic;
        prod9           : in     vl_logic;
        prod10          : in     vl_logic;
        prod11          : in     vl_logic;
        prod12          : in     vl_logic;
        prod13          : in     vl_logic;
        prod14          : in     vl_logic;
        prod15          : in     vl_logic;
        prod16          : in     vl_logic;
        prod17          : in     vl_logic;
        prod18          : in     vl_logic;
        prod19          : in     vl_logic;
        prod20          : in     vl_logic;
        prod21          : in     vl_logic;
        prod22          : in     vl_logic;
        prod23          : in     vl_logic;
        prod24          : in     vl_logic;
        prod25          : in     vl_logic;
        prod26          : in     vl_logic;
        prod27          : in     vl_logic;
        prod28          : in     vl_logic;
        prod29          : in     vl_logic;
        prod30          : in     vl_logic;
        prod31          : in     vl_logic;
        prod32          : in     vl_logic;
        prod33          : in     vl_logic;
        prod34          : in     vl_logic;
        prod35          : in     vl_logic;
        prod36          : in     vl_logic;
        prod37          : in     vl_logic;
        prod38          : in     vl_logic;
        prod39          : in     vl_logic;
        prod40          : in     vl_logic;
        prod41          : in     vl_logic;
        prod42          : in     vl_logic;
        prod43          : in     vl_logic;
        prod44          : in     vl_logic;
        prod45          : in     vl_logic;
        prod46          : in     vl_logic;
        prod47          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Multiplier_vlg_check_tst;
