library verilog;
use verilog.vl_types.all;
entity Normalizer is
    port(
        B0              : out    vl_logic;
        F0              : in     vl_logic;
        F1              : in     vl_logic;
        F2              : in     vl_logic;
        F3              : in     vl_logic;
        F4              : in     vl_logic;
        F5              : in     vl_logic;
        F6              : in     vl_logic;
        F7              : in     vl_logic;
        F8              : in     vl_logic;
        F9              : in     vl_logic;
        F10             : in     vl_logic;
        F11             : in     vl_logic;
        F12             : in     vl_logic;
        F13             : in     vl_logic;
        F14             : in     vl_logic;
        F15             : in     vl_logic;
        F16             : in     vl_logic;
        F17             : in     vl_logic;
        F18             : in     vl_logic;
        F19             : in     vl_logic;
        F20             : in     vl_logic;
        F21             : in     vl_logic;
        F22             : in     vl_logic;
        Sel             : in     vl_logic;
        Clk             : in     vl_logic;
        En              : in     vl_logic;
        F23             : in     vl_logic;
        F24             : in     vl_logic;
        F25             : in     vl_logic;
        F26             : in     vl_logic;
        F27             : in     vl_logic;
        F28             : in     vl_logic;
        F29             : in     vl_logic;
        F30             : in     vl_logic;
        F31             : in     vl_logic;
        F32             : in     vl_logic;
        F33             : in     vl_logic;
        F34             : in     vl_logic;
        F35             : in     vl_logic;
        F36             : in     vl_logic;
        F37             : in     vl_logic;
        F38             : in     vl_logic;
        F39             : in     vl_logic;
        F40             : in     vl_logic;
        F41             : in     vl_logic;
        F42             : in     vl_logic;
        F43             : in     vl_logic;
        F44             : in     vl_logic;
        F45             : in     vl_logic;
        B1              : out    vl_logic;
        B2              : out    vl_logic;
        B3              : out    vl_logic;
        B4              : out    vl_logic;
        B5              : out    vl_logic;
        B6              : out    vl_logic;
        B7              : out    vl_logic;
        B8              : out    vl_logic;
        B9              : out    vl_logic;
        B10             : out    vl_logic;
        B11             : out    vl_logic;
        B12             : out    vl_logic;
        B13             : out    vl_logic;
        B14             : out    vl_logic;
        B15             : out    vl_logic;
        B16             : out    vl_logic;
        B17             : out    vl_logic;
        B18             : out    vl_logic;
        B19             : out    vl_logic;
        B20             : out    vl_logic;
        B21             : out    vl_logic;
        Overflow        : out    vl_logic;
        Exp0            : in     vl_logic;
        Exp1            : in     vl_logic;
        Exp2            : in     vl_logic;
        Exp3            : in     vl_logic;
        Exp4            : in     vl_logic;
        Exp5            : in     vl_logic;
        Exp6            : in     vl_logic;
        Exp7            : in     vl_logic;
        E7              : out    vl_logic;
        E6              : out    vl_logic;
        E5              : out    vl_logic;
        E4              : out    vl_logic;
        E3              : out    vl_logic;
        E2              : out    vl_logic;
        E1              : out    vl_logic;
        E0              : out    vl_logic;
        B22             : out    vl_logic
    );
end Normalizer;
