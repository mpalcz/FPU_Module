library verilog;
use verilog.vl_types.all;
entity Multiplier_vlg_vec_tst is
end Multiplier_vlg_vec_tst;
